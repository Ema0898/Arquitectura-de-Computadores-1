module instruction_memory(input logic [23:0] a,
								  output logic [23:0] rd);								  
								  
<<<<<<< HEAD
  logic [23:0] memory [128];  
  
  assign memory[0] = 24'b111001101000000010001000; // MOVER R1, #8
  assign memory[1] = 24'b111001101000000010001000; // MOVER R1, #8
  assign memory[2] = 24'b111001101000000100001000; // MOVER R2, #7
  assign memory[3] = 24'b111000110000100000010000; // COMP R1, R2
  assign memory[4] = 24'b010001101000000010001010; // MOVERGT R1, #10
  assign memory[5] = 24'b111000000000100000010000; // SUM R0, R1, R2
=======
  logic [23:0] memory [140];
	/*initial
		$readmemb("instructions.dat", memory);  */
  
  /*assign memory[0] = 24'b111001101000000010001000; // MOVER R1, #8
  assign memory[1] = 24'b111001101000000010001000; // MOVER R1, #9
  assign memory[2] = 24'b111001101000000100001000; // MOVER R2, #8
  assign memory[3] = 24'b111001101000001000000010; // MOVER R4, #1
  assign memory[4] = 24'b111011111010001010000000; // LOAD R5, [R4]
  assign memory[5] = 24'b111001001010101010000001; // MUL R5, R5, 1
  assign memory[6] = 24'b111000111010100000000000; // COMP R1, 0
  assign memory[7] = 24'b001001101000000010001010; // MOVNEG R1, #10  
  assign memory[8] = 24'b111000000000100000010000; // SUM R0, R1, R2*/
>>>>>>> c9ba90840e60ad14c5f5ff539c15feeba067e3e4
  
  /*assign memory[0] = 22'b1001101000000010001000; // MOVER R1, #8
  assign memory[1] = 22'b1001101000000010001000; // MOVER R1, #8
  assign memory[2] = 22'b1001101000000100001001; // MOVER R2, #9
  assign memory[3] = 22'b1000000000100000010000; // SUM R0, R1, R2
  assign memory[4] = 22'b1011100000100000010000; // STORE R0, [R1, R2]
  assign memory[5] = 22'b1011101000100000000111; // STORE R0, [R1, #7]
  assign memory[6] = 22'b1011110000100110010000; // LOAD R3, [R1, R2]
  assign memory[7] = 22'b1011111000101000000111; // LOAD R4, [R1, #7]
  assign memory[8] = 22'b1000000001101010100000; // SUM R5, R4, R3  
  assign memory[9] = 22'b1000001010101010001111; // SUM R5, R5, #15
  assign memory[10] = 22'b1001000010101100001000;  // MUL R6, R5, R1
  assign memory[11] = 22'b1001001010001110000011; //MUL R7, R4, #3
  assign memory[12] = 22'b1000111011100000110010; // CMP R7, #50
  assign memory[13] = 22'b1001101000010000000000; // MOVER R8, #0
  assign memory[14] = 22'b0000001011110000000010; // SUMIG R8, R7, #2 // Si se ejecuta
  assign memory[15] = 22'b1000001100010000000001; // SUM R8, R8, #1*/
  
  /*assign memory[0] = 24'b111001101000000010001000; // MOVER R1, #8
  assign memory[1] = 24'b111001101000000010001000; // MOVER R1, #8
  assign memory[2] = 24'b111001101000000100001001; // MOVER R2, #9
  assign memory[3] = 24'b111001101000000110000001; // MOVER R3, #50
  assign memory[4] = 24'b111001101000001000000010; // MOVER R4, #60
  assign memory[5] = 24'b111011111001101010000000; // LOAD R5, [R3]
  assign memory[6] = 24'b111011111010001100000000; // LOAD R6, [R4]*/
  
  
  /*assign memory[0] = 24'b111001101000000110000000; // MOVER R3, #0 : Init
  assign memory[1] = 24'b111001101000000010000001; // MOVER R1, #0
  assign memory[2] = 24'b111001101000000100000001; // MOVER R2, #1
  assign memory[3] = 24'b111000110000100000010000; // COMP R1, R2
  assign memory[4] = 24'b000101111111111111101000; // SALTOIG Init
  assign memory[5] = 24'b111000001000100010000100; // SUM R1, R1, #4
  assign memory[6] = 24'b111000001001000100000101; // SUM R2, R2, #5 : Hola
  assign memory[7] = 24'b111000001000100010000111; // SUM R1, R1, #7 : Adios*/
  
  // VGA primera prueba  
  /*assign memory[0] = 22'b1001101000000000000000;
  assign memory[1] = 22'b1001101000000000000000;
  assign memory[2] = 22'b1001101000000011110100;
  assign memory[3] = 22'b1011101000100000000000;
  assign memory[4] = 22'b1001101000000001101110;
  assign memory[5] = 22'b1011111000000010000000;
  assign memory[6] = 22'b1000111000100000000001;
  assign memory[7] = 22'b0100000000000000000000;
  assign memory[8] = 22'b1101111111111111101000;
  assign memory[9] = 22'b1001101000000000000001;
  assign memory[10] = 22'b1001101000000011110100;
  assign memory[11] = 22'b1011101000100000000000;
  assign memory[12] = 22'b1101111111111111011000;*/
  
  
  // Ultima prueba simulacion
  /*assign memory[0] = 22'b01001101000000000000000;
  assign memory[1] = 22'b01001101000000000000000;
  assign memory[2] = 22'b1001101000000011110100;
  assign memory[3] = 22'b1011101000100000000000;
  assign memory[4] = 22'b1001101000000000000001;
  assign memory[5] = 22'b1001101000000011111001;
  assign memory[6] = 22'b1011101000100000000000;
  assign memory[7] = 22'b1001101000000111101000;
  assign memory[8] = 22'b1011111000100000000000;
  assign memory[9] = 22'b1011111001100100000000;
  assign memory[10] = 22'b1000110001000000000000;
  assign memory[11] = 22'b0100000000000000000000;
  assign memory[12] = 22'b1101111111111111100100;
  assign memory[13] = 22'b1001101000000000000001;
  assign memory[14] = 22'b1001101000000101110100;
  assign memory[15] = 22'b1011101001000000000000;
  assign memory[16] = 22'b1101111111111111010100;*/
  
  // Ultima prueba  
  /*assign memory[0] = 22'b1001101000000000000000;
  assign memory[1] = 22'b1001101000000000000000;
  assign memory[2] = 22'b1001101000000011110100;
  assign memory[3] = 22'b1011101000100000000000;
  assign memory[4] = 22'b1001101000000000000001;
  assign memory[5] = 22'b1001101000000011111001;
  assign memory[6] = 22'b1011101000100000000000;
  assign memory[7] = 22'b1011111000100000000000;
  assign memory[8] = 22'b1000111000000000000001;
  assign memory[9] = 22'b0100000000000000000000;
  assign memory[10] = 22'b1101111111111111101100;
  assign memory[11] = 22'b1001101000000000000001;
  assign memory[12] = 22'b1001101000000101110100;
  assign memory[13] = 22'b1011101001000000000000;
  assign memory[14] = 22'b1101111111111111011100;*/
 
  
  // Prueba boton leyendo de memoria  
  /*assign memory[0] = 22'b1001101000000000000000;
  assign memory[1] = 22'b1001101000000000000000;
  assign memory[2] = 22'b1001101000000011110100;
  assign memory[3] = 22'b1011101000100000000000;
  assign memory[4] = 22'b1001101000000000000001;
  assign memory[5] = 22'b1001101000000011111001;
  assign memory[6] = 22'b1011101000100000000000;
  assign memory[7] = 22'b1001101000000111101000;
  assign memory[8] = 22'b1011111000100000000000;
  assign memory[9] = 22'b1011111001100100000000;
  assign memory[10] = 22'b1000110001000000000000;
  assign memory[11] = 22'b0100000000000000000000;
  assign memory[12] = 22'b1101111111111111100100;
  assign memory[13] = 22'b1001101000000000000001;
  assign memory[14] = 22'b1001101000000101110100;
  assign memory[15] = 22'b1011101001000000000000;
  assign memory[16] = 22'b1101111111111111010100;*/
  
  // Prueba boton leyendo de memoria 2
  
  /*assign memory[0] = 22'b1001101000000000000000;
  assign memory[1] = 22'b1001101000000000000000;
  assign memory[2] = 22'b1001101000000011110100;
  assign memory[3] = 22'b1011101000100000000000;
  assign memory[4] = 22'b1001101000000000000001;
  assign memory[5] = 22'b1001101000000011010011;
  assign memory[6] = 22'b1001001000100010110010;
  assign memory[7] = 22'b1001101000000100101000;
  assign memory[8] = 22'b1001001001000100000011;
  assign memory[9] = 22'b1000000000100010010000;
  assign memory[10] = 22'b1011101000100000000000;
  assign memory[11] = 22'b1001101000000111101000;
  assign memory[12] = 22'b1011111000100000000000;
  assign memory[13] = 22'b1011111001100100000000;
  assign memory[14] = 22'b1000110001000000000000;
  assign memory[15] = 22'b0100000000000000000000;
  assign memory[16] = 22'b1101111111111111100100;
  assign memory[17] = 22'b1001101000000000000001;
  assign memory[18] = 22'b1001101000000101110100;
  assign memory[19] = 22'b1011101001000000000000;
  assign memory[20] = 22'b1101111111111111010100;*/
  
  assign memory[0] = 24'b111001101000000100000000;
	assign memory[1] = 24'b111001101000000100000000;
	assign memory[2] = 24'b111001101000000011101000;
	assign memory[3] = 24'b111011111000100000000000;
	assign memory[4] = 24'b111000111000000000000001;
	assign memory[5] = 24'b000100000000000000101000;
	assign memory[6] = 24'b111000001001000100001001;
	assign memory[7] = 24'b111000001000100010000100;
	assign memory[8] = 24'b111011111000100000000000;
	assign memory[9] = 24'b111000111000000000000001;
	assign memory[10] = 24'b000100000000000000010100;
	assign memory[11] = 24'b111000001001000100001001;
	assign memory[12] = 24'b111000001000100010000100;
	assign memory[13] = 24'b111011111000100000000000;
	assign memory[14] = 24'b111000111000000000000001;
	assign memory[15] = 24'b000100000000000000000000;
	assign memory[16] = 24'b111101111111111110111000;
	assign memory[17] = 24'b111001101000000001110100;
	assign memory[18] = 24'b111001101000000010000000;
	assign memory[19] = 24'b111011101000000010000000;
	assign memory[20] = 24'b111001101000001011111111;
	assign memory[21] = 24'b111001101000000000000000;
	assign memory[22] = 24'b111001101000000011100100;
	assign memory[23] = 24'b111000001000100011100100;
	assign memory[24] = 24'b111000001000100011100100;
	assign memory[25] = 24'b111000001000100011100100;
	assign memory[26] = 24'b111001101000000111111000;
	assign memory[27] = 24'b111001101000001001010000;
	assign memory[28] = 24'b111001001010001000110010;
	assign memory[29] = 24'b111000001010001000000011;
	assign memory[30] = 24'b111001001010001000101000;
	assign memory[31] = 24'b111101111111111111111100;
	assign memory[32] = 24'b111000110000000000001000;
	assign memory[33] = 24'b000100000000000000010100;
	assign memory[34] = 24'b111011101010001010000000;
	assign memory[35] = 24'b111000001010001000000001;
	assign memory[36] = 24'b111000001000000000000001;
	assign memory[37] = 24'b111001101000001100000000;
	assign memory[38] = 24'b111001101000001110000010;
	assign memory[39] = 24'b111101111111111111011100;
	assign memory[40] = 24'b111001101000000011100100;
	assign memory[41] = 24'b111000001000100011100100;
	assign memory[42] = 24'b111000001000100011100100;
	assign memory[43] = 24'b111000001000100011100100;
	assign memory[44] = 24'b111001101000001011111111;
	assign memory[45] = 24'b111000110011100000001000;
	assign memory[46] = 24'b000100000000000000010000;
	assign memory[47] = 24'b111000110011000000001000;
	assign memory[48] = 24'b000100000000000000110100;
	assign memory[49] = 24'b111000111011000000000000;
	assign memory[50] = 24'b000100000000000001000100;
	assign memory[51] = 24'b111100000000000001010000;
	assign memory[52] = 24'b111001101000000000000000;
	assign memory[53] = 24'b111000110000000000001000;
	assign memory[54] = 24'b000100000000000000001100;
	assign memory[55] = 24'b111011101010001010000000;
	assign memory[56] = 24'b111000001010001000000001;
	assign memory[57] = 24'b111000001000000000000001;
	assign memory[58] = 24'b111101111111111111100100;
	assign memory[59] = 24'b111001101000000001110100;
	assign memory[60] = 24'b111001101000000010000001;
	assign memory[61] = 24'b111011101000000010000000;
	assign memory[62] = 24'b111101111111111100000000;
	assign memory[63] = 24'b111011101010001010000000;
	assign memory[64] = 24'b111000001010001000000001;
	assign memory[65] = 24'b111000001011101110000001;
	assign memory[66] = 24'b111000001001100110000010;
	assign memory[67] = 24'b111001101000001100000000;
	assign memory[68] = 24'b111101111111111110011100;
	assign memory[69] = 24'b111011101010001010000000;
	assign memory[70] = 24'b111000001010001000000001;
	assign memory[71] = 24'b111000001011001100000010;
	assign memory[72] = 24'b111101111111111110001100;
	assign memory[73] = 24'b111001101000000010000000;
	assign memory[74] = 24'b111001101000001010000000;
	assign memory[75] = 24'b111011111001000000000000;
	assign memory[76] = 24'b111011111001110010000000;
	assign memory[77] = 24'b111001000000010101001000;
	assign memory[78] = 24'b111000000000100011010000;
	assign memory[79] = 24'b111000001010101010000001;
	assign memory[80] = 24'b111011111001000000000001;
	assign memory[81] = 24'b111011110001110010101000;
	assign memory[82] = 24'b111001000000010101001000;
	assign memory[83] = 24'b111000000000100011010000;
	assign memory[84] = 24'b111000001010101010000001;
	assign memory[85] = 24'b111011111001000000000010;
	assign memory[86] = 24'b111011110001110010101000;
	assign memory[87] = 24'b111001000000010101001000;
	assign memory[88] = 24'b111000000000100011010000;
	assign memory[89] = 24'b111000001010101011100100;
	assign memory[90] = 24'b111000001010101011100100;
	assign memory[91] = 24'b111000001010101011100100;
	assign memory[92] = 24'b111000001010101011100010;
	assign memory[93] = 24'b111011111001000000000011;
	assign memory[94] = 24'b111011110001110010101000;
	assign memory[95] = 24'b111001000000010101001000;
	assign memory[96] = 24'b111000000000100011010000;
	assign memory[97] = 24'b111000001010101010000001;
	assign memory[98] = 24'b111011111001000000000100;
	assign memory[99] = 24'b111011110001110010101000;
	assign memory[100] = 24'b111001000000010101001000;
	assign memory[101] = 24'b111000000000100011010000;
	assign memory[102] = 24'b111000001010101010000001;
	assign memory[103] = 24'b111011111001000000000101;
	assign memory[104] = 24'b111011110001110010101000;
	assign memory[105] = 24'b111001000000010101001000;
	assign memory[106] = 24'b111000000000100011010000;
	assign memory[107] = 24'b111000001010101011100100;
	assign memory[108] = 24'b111000001010101011100100;
	assign memory[109] = 24'b111000001010101011100100;
	assign memory[110] = 24'b111000001010101011100010;
	assign memory[111] = 24'b111011111001000000000110;
	assign memory[112] = 24'b111011110001110010101000;
	assign memory[113] = 24'b111001000000010101001000;
	assign memory[114] = 24'b111000000000100011010000;
	assign memory[115] = 24'b111000001010101010000001;
	assign memory[116] = 24'b111011111001000000000111;
	assign memory[117] = 24'b111011110001110010101000;
	assign memory[118] = 24'b111001000000010101001000;
	assign memory[119] = 24'b111000000000100011010000;
	assign memory[120] = 24'b111000001010101010000001;
	assign memory[121] = 24'b111011111001000000001000;
	assign memory[122] = 24'b111011110001110010101000;
	assign memory[123] = 24'b111001000000010101001000;
	assign memory[124] = 24'b111000000000100011010000;
	assign memory[125] = 24'b111001101000010000000000;
	assign memory[126] = 24'b111000110000100001000000;
	assign memory[127] = 24'b001001101000000010000000;
	assign memory[128] = 24'b111000001100010001100100;
	assign memory[129] = 24'b111000001100010001100100;
	assign memory[130] = 24'b111000001100010000110111;
	assign memory[131] = 24'b111000110000100001000000;
	assign memory[132] = 24'b010001101000000011100100;
	assign memory[133] = 24'b010000001000100011100100;
	assign memory[134] = 24'b010000001000100010110111;
	assign memory[135] = 24'b111011101010000010000000;
	assign memory[136] = 24'b111000001001100110000001;
	assign memory[137] = 24'b111000001010001000000001;
	assign memory[138] = 24'b111000001011001100000001;
	assign memory[139] = 24'b111101111111111001101100;
	
  assign rd = memory[a[21:2]]; // word aligned
			  
endmodule 
