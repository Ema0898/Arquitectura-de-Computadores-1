module decode_unit(input logic cond,
						input logic [1:0] op,
						input logic [2:0] funct,
						input logic [3:0] rd,
						output logic pc_src, reg_write, mem_write, mem_reg, alu_src, no_write, mov_src, reg_src,
						output logic [1:0] alu_control, imm_src, flag_write);

	

endmodule 